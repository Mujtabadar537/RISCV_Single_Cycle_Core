module AND_Gate(

input in1_i,
input in2_i,

output  out_o

);


assign out_o = in1_i & in2_i;


endmodule
